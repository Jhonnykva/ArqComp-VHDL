library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port( clk : in std_logic;
        endereco : in unsigned(6 downto 0);--memória de programa = 4Kbytes 4000bytes = 32000 bits
        instr : out unsigned(16 downto 0)    --32000/17=1882 endereços de 17 bits
    );
end entity;

architecture a_rom of rom is
    type mem is array (0 to 127) of unsigned(16 downto 0);--trocar futuramente 127 por 1881
    constant conteudo_rom : mem := (
        -- caso endereco => conteudo
        0 => B"00001100_000000001",
        1 => B"01001_011_000000001",
        2 => B"00000011_000000011",
        3 => B"00001010_000000000",
        4 => B"00001101_000000000",
        5 => B"00001110_000000001",
        6 => B"00000010_000000011",
        7 => B"00000111_000000000",
        8 => B"00000101_000100001",
        9 => B"00001000_011111000",
        10=> B"00001100_000000100",
        11=> B"01001_011_000000100",
        12=> B"00000001_000000000",
        13=> B"00001010_000000000",
        14=> B"00001101_000000000",
        15=> B"00001101_000000000",
        16=> B"00000011_000000011",
        17=> B"00001110_000000010",
        18=> B"00000010_000000011",
        19=> B"00000111_000000000",
        20=> B"00000101_000100001",
        21=> B"00001000_011110110",
        22=> B"00001100_000000110",
        23=> B"01001_011_000000110",
        24=> B"00000001_000000000",
        25=> B"00001010_000000000",
        26=> B"00001101_000000000",
        27=> B"00001101_000000000",
        28=> B"00001101_000000000",
        29=> B"00000011_000000011",
        30=> B"00001110_000000011",
        31=> B"00000010_000000011",
        32=> B"00000111_000000000",
        33=> B"00000101_000100001",
        34=> B"00001000_011110101",
        35=> B"00001100_000001010",
        36=> B"01001_011_000001010",
        37=> B"00000001_000000000",
        38=> B"00001010_000000000",
        39=> B"00001101_000000000",
        40=> B"00001101_000000000",
        41=> B"00001101_000000000",
        42=> B"00001101_000000000",
        43=> B"00001101_000000000",
        44=> B"00000011_000000011",
        45=> B"00001110_000000101",
        46=> B"00000010_000000011",
        47=> B"00000111_000000000",
        48=> B"00000101_000100001",
        49=> B"00001000_011110011",
        50=> B"00001100_000000010",
        51=> B"01001_100_000000010",
        52=> B"00001011_000000000",
        53=> B"00000010_000000101",
        54=> B"00000011_000000100",
        55=> B"00001110_000000001",
        56=> B"00001101_000000000",
        57=> B"00000010_000000100",
        58=> B"00000111_000000000",
        59=> B"00000101_000100001",
        60=> B"00001000_011110111",
        -- abaixo: casos omissos => (zero em todos os bits)
        others => (others=>'0')
    );

begin
    process(clk)
    begin
        if(rising_edge(clk)) then
        instr <= conteudo_rom(to_integer(endereco));
    end if;
end process;
end architecture;