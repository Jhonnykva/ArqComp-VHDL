$date
  Wed Nov 03 22:23:54 2021
$end
$version
  GHDL v0
$end
$timescale
  1 fs
$end
$scope module standard $end
$upscope $end
$scope module std_logic_1164 $end
$upscope $end
$scope module numeric_std $end
$upscope $end
$scope module gerenciador_tb $end
$var reg 16 ! reg_in_1[15:0] $end
$var reg 16 " reg_in_2[15:0] $end
$var reg 16 # reg_out[15:0] $end
$var reg 3 $ select_reg_1[2:0] $end
$var reg 3 % select_reg_2[2:0] $end
$var reg 3 & select_reg_3[2:0] $end
$var reg 1 ' rst_reg $end
$scope module uut $end
$var reg 16 ( reg_in_1[15:0] $end
$var reg 16 ) reg_in_2[15:0] $end
$var reg 16 * reg_out[15:0] $end
$var reg 3 + select_reg_1[2:0] $end
$var reg 3 , select_reg_2[2:0] $end
$var reg 3 - select_reg_3[2:0] $end
$var reg 1 . rst_reg $end
$var reg 1 / finished $end
$var reg 1 0 clk $end
$var reg 1 1 reset $end
$var reg 1 2 wr_enable_1 $end
$var reg 1 3 wr_enable_2 $end
$var reg 1 4 wr_enable_3 $end
$var reg 1 5 wr_enable_4 $end
$var reg 1 6 wr_enable_5 $end
$var reg 1 7 wr_enable_6 $end
$var reg 1 8 wr_enable_7 $end
$var reg 1 9 wr_enable_0 $end
$var reg 16 : data_in_1[15:0] $end
$var reg 16 ; data_in_2[15:0] $end
$var reg 16 < data_in_3[15:0] $end
$var reg 16 = data_in_4[15:0] $end
$var reg 16 > data_in_5[15:0] $end
$var reg 16 ? data_in_6[15:0] $end
$var reg 16 @ data_in_7[15:0] $end
$var reg 16 A data_out_1[15:0] $end
$var reg 16 B data_out_2[15:0] $end
$var reg 16 C data_out_3[15:0] $end
$var reg 16 D data_out_4[15:0] $end
$var reg 16 E data_out_5[15:0] $end
$var reg 16 F data_out_6[15:0] $end
$var reg 16 G data_out_7[15:0] $end
$var reg 16 H data_out_0[15:0] $end
$scope module reg1 $end
$var reg 1 I clk $end
$var reg 1 J rst $end
$var reg 1 K wr_enable $end
$var reg 16 L data_in[15:0] $end
$var reg 16 M data_out[15:0] $end
$var reg 16 N registro[15:0] $end
$upscope $end
$scope module reg2 $end
$var reg 1 O clk $end
$var reg 1 P rst $end
$var reg 1 Q wr_enable $end
$var reg 16 R data_in[15:0] $end
$var reg 16 S data_out[15:0] $end
$var reg 16 T registro[15:0] $end
$upscope $end
$scope module reg3 $end
$var reg 1 U clk $end
$var reg 1 V rst $end
$var reg 1 W wr_enable $end
$var reg 16 X data_in[15:0] $end
$var reg 16 Y data_out[15:0] $end
$var reg 16 Z registro[15:0] $end
$upscope $end
$scope module reg4 $end
$var reg 1 [ clk $end
$var reg 1 \ rst $end
$var reg 1 ] wr_enable $end
$var reg 16 ^ data_in[15:0] $end
$var reg 16 _ data_out[15:0] $end
$var reg 16 ` registro[15:0] $end
$upscope $end
$scope module reg5 $end
$var reg 1 a clk $end
$var reg 1 b rst $end
$var reg 1 c wr_enable $end
$var reg 16 d data_in[15:0] $end
$var reg 16 e data_out[15:0] $end
$var reg 16 f registro[15:0] $end
$upscope $end
$scope module reg6 $end
$var reg 1 g clk $end
$var reg 1 h rst $end
$var reg 1 i wr_enable $end
$var reg 16 j data_in[15:0] $end
$var reg 16 k data_out[15:0] $end
$var reg 16 l registro[15:0] $end
$upscope $end
$scope module reg7 $end
$var reg 1 m clk $end
$var reg 1 n rst $end
$var reg 1 o wr_enable $end
$var reg 16 p data_in[15:0] $end
$var reg 16 q data_out[15:0] $end
$var reg 16 r registro[15:0] $end
$upscope $end
$scope module reg0 $end
$var reg 1 s clk $end
$var reg 1 t rst $end
$var reg 1 u wr_enable $end
$var reg 16 v data_in[15:0] $end
$var reg 16 w data_out[15:0] $end
$var reg 16 x registro[15:0] $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
bUUUUUUUUUUUUUUUU !
bUUUUUUUUUUUUUUUU "
b0000000000001110 #
bUUU $
bUUU %
b110 &
U'
bUUUUUUUUUUUUUUUU (
bUUUUUUUUUUUUUUUU )
b0000000000001110 *
bUUU +
bUUU ,
b110 -
U.
0/
U0
U1
02
03
04
05
06
17
08
09
bUUUUUUUUUUUUUUUU :
bUUUUUUUUUUUUUUUU ;
bUUUUUUUUUUUUUUUU <
bUUUUUUUUUUUUUUUU =
bUUUUUUUUUUUUUUUU >
bUUUUUUUUUUUUUUUU ?
bUUUUUUUUUUUUUUUU @
bUUUUUUUUUUUUUUUU A
bUUUUUUUUUUUUUUUU B
bUUUUUUUUUUUUUUUU C
bUUUUUUUUUUUUUUUU D
bUUUUUUUUUUUUUUUU E
bUUUUUUUUUUUUUUUU F
bUUUUUUUUUUUUUUUU G
bUUUUUUUUUUUUUUUU H
UI
UJ
0K
bUUUUUUUUUUUUUUUU L
bUUUUUUUUUUUUUUUU M
bUUUUUUUUUUUUUUUU N
UO
UP
0Q
bUUUUUUUUUUUUUUUU R
bUUUUUUUUUUUUUUUU S
bUUUUUUUUUUUUUUUU T
UU
UV
0W
bUUUUUUUUUUUUUUUU X
bUUUUUUUUUUUUUUUU Y
bUUUUUUUUUUUUUUUU Z
U[
U\
0]
bUUUUUUUUUUUUUUUU ^
bUUUUUUUUUUUUUUUU _
bUUUUUUUUUUUUUUUU `
Ua
Ub
0c
bUUUUUUUUUUUUUUUU d
bUUUUUUUUUUUUUUUU e
bUUUUUUUUUUUUUUUU f
Ug
Uh
1i
bUUUUUUUUUUUUUUUU j
bUUUUUUUUUUUUUUUU k
bUUUUUUUUUUUUUUUU l
Um
Un
0o
bUUUUUUUUUUUUUUUU p
bUUUUUUUUUUUUUUUU q
bUUUUUUUUUUUUUUUU r
Us
Ut
0u
b0000000000000000 v
bUUUUUUUUUUUUUUUU w
bUUUUUUUUUUUUUUUU x
#50000000
b0000000000000000 #
b100 &
b0000000000000000 *
b100 -
15
07
1]
0i
#100000000
b0000000000001110 #
b110 &
b0000000000001110 *
b110 -
05
17
0]
1i
#150000000
b0000000000000000 #
b100 &
b0000000000000000 *
b100 -
15
07
1]
0i
#200000000
